module WB_Stage(output out);
  assign out = 1;
endmodule
