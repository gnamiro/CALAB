module ConditionCheck(
  input [3:0] cond, Sr,
  output condRes
);

assign condRes = 1'b0;

endmodule
